module rca_nbit #(
	parameter N = 64
)(
	input		[N-1:0] i_a,
	input		[N-1:0] i_b,
	input				i_c,
	output wire [N-1:0] o_s,
	output wire			o_c
);

	wire [N-1:0] p;
	wire [N-1:0] g;
	// verilator lint_off UNOPTFLAT
	wire [N:0] c;
	// verilator lint_on UNOPTFLAT

	genvar i;
	for (i = 0; i < N; i = i+1) begin: csa
		assign g[i]   = i_a[i] & i_b[i];
		assign p[i]   = i_a[i] ^ i_b[i];
		assign c[i+1] = c[i] & p[i] | g[i];
		assign o_s[i] = p[i] ^ c[i];
	end

	assign c[0] = i_c;
	assign o_c = c[N];

endmodule